*
*
*
*                       LINUX           Fri Oct 24 13:35:10 2025
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 24.1.0-p089
*  Build Date     : Wed Dec 18 09:06:09 PST 2024
*
*  HSPICE LIBRARY
*
*  QRC_TECH_DIR /ece558_658/pdk/verification/qrc/typical 
*
*
*

*
.SUBCKT XOR_X1 CIN COUT GND PHI RST SOUT VDD
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MNM23	net1#14	net7#3	net12#4	GND	g45n1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM13	net2#21	CIN#6	net37#3	GND	g45n1svt
+ L=4.5e-08	W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM26	net21#4	net1#3	GND#20	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM14	net33#4	net6#2	GND#13	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM25	net8#5	PHI#6	net21#2	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM21	net10#4	RST#1	GND#10	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM12	net2#6	net3#3	net33#2	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM24	net12	net4#3	GND#7	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM15	net37	SOUT#3	GND#6	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM20	net4#5	net2	net10#2	GND	g45n1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.52678 scb=0.000111658 scc=3.66286e-09 fw=2.4e-07
MNM27	net7#7	PHI#3	GND#2	GND	g45n1svt	L=4.5e-08
+ W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=5.20631 scb=0.0011851 scc=1.90632e-06 fw=1.2e-07
MNM10	net3#8	CIN#1	GND#3	GND	g45n1svt	L=4.5e-08
+ W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MNM11	net6#6	SOUT#4	GND#12	GND	g45n1svt	L=4.5e-08
+ W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MNM28	COUT#2	net6#4	GND#15	GND	g45n1svt	L=4.5e-08
+ W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MNM22	SOUT#10	net8	GND#18	GND	g45n1svt	L=4.5e-08
+ W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MNM29	COUT#8	net3#4	GND#21	GND	g45n1svt	L=4.5e-08
+ W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
+ sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 fw=1.2e-07
MPM25	net7#4	PHI#1	VDD#2	VDD	g45p1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=6.96428 scb=0.00265505 scc=6.98372e-06 fw=2.4e-07
MPM10	net3#10	CIN#3	VDD#4	VDD	g45p1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=11.4009 scb=0.010956 scc=0.000489739 fw=2.4e-07
MPM18	net4#6	net2#3	VDD#5	VDD	g45p1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.05637 scb=0.0041121 scc=4.83436e-05 fw=2.4e-07
MPM13	net13#6	SOUT#1	VDD#9	VDD	g45p1svt	L=4.5e-08
+ W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=6.03189 scb=0.00286778 scc=3.79924e-05 fw=4.8e-07
MPM22	net27#6	net4	VDD#14	VDD	g45p1svt	L=4.5e-08
+ W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=6.25222 scb=0.0032094 scc=4.93602e-05 fw=4.8e-07
MPM14	net2#10	net3	net13#3	VDD	g45p1svt
+ L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=6.03189 scb=0.00286778 scc=3.79924e-05 fw=4.8e-07
MPM19	net4#10	RST#3	VDD#18	VDD	g45p1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=7.05637 scb=0.0041121 scc=4.83436e-05 fw=2.4e-07
MPM11	net6#8	SOUT#6	VDD#19	VDD	g45p1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=11.971 scb=0.0117186 scc=0.000577399 fw=2.4e-07
MPM21	net1#6	PHI#4	net27#3	VDD	g45p1svt	L=4.5e-08
+ W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=6.25222 scb=0.0032094 scc=4.93602e-05 fw=4.8e-07
MPM29	COUT#5	net6#5	net14#3	VDD	g45p1svt	L=4.5e-08
+ W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=7.78706 scb=0.00554847 scc=0.000178111 fw=4.8e-07
MPM12	net18#3	net6	VDD#23	VDD	g45p1svt	L=4.5e-08
+ W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=6.03189 scb=0.00286778 scc=3.79924e-05 fw=4.8e-07
MPM20	SOUT#12	net8#3	VDD#27	VDD	g45p1svt	L=4.5e-08
+ W=2.4e-07
+ AD=3.36e-14	AS=3.36e-14	PD=7.6e-07	PS=7.6e-07
+ sa=1.4e-07 sb=1.4e-07 sca=11.6789 scb=0.0113323 scc=0.000531848 fw=2.4e-07
MPM23	net5#5	net1	VDD#30	VDD	g45p1svt	L=4.5e-08
+ W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=6.4958 scb=0.00358872 scc=6.40322e-05 fw=4.8e-07
MPM28	net14#7	net3#6	VDD#35	VDD	g45p1svt	L=4.5e-08
+ W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=7.52782 scb=0.0051674 scc=0.00015053 fw=4.8e-07
MPM15	net2#15	CIN#4	net18#8	VDD	g45p1svt
+ L=4.5e-08	W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=6.03189 scb=0.00286778 scc=3.79924e-05 fw=4.8e-07
MPM24	net8#10	net7	net5#3	VDD	g45p1svt	L=4.5e-08
+ W=4.8e-07
+ AD=6.72e-14	AS=6.72e-14	PD=1.24e-06	PS=1.24e-06
+ sa=1.4e-07 sb=1.4e-07 sca=7.06783 scb=0.00447348 scc=0.000107211 fw=4.8e-07
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rl1	PHI#1	PHI#2	285.713379	$poly_conn
Rl2	PHI#2	PHI#3	62.636475	$poly_conn
Rl3	CIN#1	CIN#2	167.287628	$poly_conn
Rl4	CIN#2	CIN#3	236.518387	$poly_conn
Rl5	net2	net2#2	53.021091	$poly_conn
Rl6	net2#2	net2#3	272.251862	$poly_conn
Rl7	SOUT#1	SOUT#2	211.518387	$poly_conn
Rl8	SOUT#2	SOUT#3	67.287621	$poly_conn
Rl9	net4	net4#2	53.826080	$poly_conn
Rl10	net4#2	net4#3	207.672241	$poly_conn
Rl11	net3	net3#2	126.098015	$poly_conn
Rl12	net3#2	net3#3	151.098022	$poly_conn
Rl13	RST#1	RST#2	161.518402	$poly_conn
Rl14	RST#2	RST#3	165.364548	$poly_conn
Rl15	SOUT#4	SOUT#5	339.559540	$poly_conn
Rl16	SOUT#5	SOUT#6	58.790321	$poly_conn
Rl17	PHI#4	PHI#5	221.133774	$poly_conn
Rl18	PHI#5	PHI#6	63.441463	$poly_conn
Rl19	net6	net6#2	340.384613	$poly_conn
Rl20	net6#2	net6#3	376.902985	$poly_conn
Rl21	net6#3	net6#4	138.441452	$poly_conn
Rl22	net6#4	net6#5	303.846161	$poly_conn
Rl23	net8	net8#2	242.287628	$poly_conn
Rl24	net8#2	net8#3	159.595306	$poly_conn
Rl25	net1	net1#2	55.749157	$poly_conn
Rl26	net1#2	net1#3	219.210693	$poly_conn
Rl27	net3#4	net3#5	215.364548	$poly_conn
Rl28	net3#5	net3#6	53.826077	$poly_conn
Rl29	CIN#4	CIN#5	209.595322	$poly_conn
Rl30	CIN#5	CIN#6	69.210693	$poly_conn
Rl31	net7	net7#2	134.595322	$poly_conn
Rl32	net7#2	net7#3	128.826080	$poly_conn
Rk1	VDD#1	VDD#2	31.001551	$metal1_conn
Rk2	GND#1	GND#2	75.002892	$metal1_conn
Rk3	net7#4	net7#5	31.000000	$metal1_conn
Rk4	net7#6	net7#7	75.002892	$metal1_conn
Rk5	GND#3	GND#4	75.000000	$metal1_conn
Rk6	VDD#3	VDD#4	31.004650	$metal1_conn
Rk7	net10	net10#2	37.501549	$metal1_conn
Rk8	VDD#5	VDD#6	31.000000	$metal1_conn
Rk9	VDD#7	VDD#8	0.160332	$metal1_conn
Rk10	VDD#8	VDD#10	0.009138	$metal1_conn
Rk11	VDD#10	VDD#11	0.173343	$metal1_conn
Rk12	VDD#9	VDD#10	15.500000	$metal1_conn
Rk13	GND#5	GND#6	37.501549	$metal1_conn
Rk14	net3#7	net3#8	75.002892	$metal1_conn
Rk15	net3#9	net3#10	31.004650	$metal1_conn
Rk16	net2#2	net2#5	45.306679	$metal1_conn
Rk17	SOUT#2	SOUT#8	45.521744	$metal1_conn
Rk18	net4#4	net4#5	37.501549	$metal1_conn
Rk19	net4#6	net4#7	31.000000	$metal1_conn
Rk20	net37	net37#2	37.500000	$metal1_conn
Rk21	GND#7	GND#8	37.511574	$metal1_conn
Rk22	VDD#12	VDD#13	0.160250	$metal1_conn
Rk23	VDD#13	VDD#15	0.002894	$metal1_conn
Rk24	VDD#15	VDD#16	0.164837	$metal1_conn
Rk25	VDD#14	VDD#15	15.500000	$metal1_conn
Rk26	net12	net12#2	37.511574	$metal1_conn
Rk27	net4#2	net4#9	45.249928	$metal1_conn
Rk28	net33	net33#2	37.501549	$metal1_conn
Rk29	net13	net13#2	0.153140	$metal1_conn
Rk30	net13#2	net13#4	0.003215	$metal1_conn
Rk31	net13#4	net13#5	0.652994	$metal1_conn
Rk32	net13#5	net13#7	0.001039	$metal1_conn
Rk33	net13#7	net13#8	0.153858	$metal1_conn
Rk34	net13#4	net13#9	0.156763	$metal1_conn
Rk35	net13#3	net13#4	15.500000	$metal1_conn
Rk36	net13#6	net13#7	15.500000	$metal1_conn
Rk37	GND#9	GND#10	37.503101	$metal1_conn
Rk38	VDD#17	VDD#18	31.001551	$metal1_conn
Rk39	RST#2	RST	46.321747	$metal1_conn
Rk40	GND#11	GND#12	75.002892	$metal1_conn
Rk41	VDD#19	VDD#20	31.001551	$metal1_conn
Rk42	net2#6	net2#7	37.500000	$metal1_conn
Rk43	net2#8	net2#9	0.160250	$metal1_conn
Rk44	net2#9	net2#11	0.002894	$metal1_conn
Rk45	net2#11	net2#12	0.164837	$metal1_conn
Rk46	net2#10	net2#11	15.500000	$metal1_conn
Rk47	net10#3	net10#4	37.501549	$metal1_conn
Rk48	net4#10	net4#11	31.000000	$metal1_conn
Rk49	net10#5	net10#6	1.096976	$metal1_conn
Rk50	net4#12	net4#13	0.459784	$metal1_conn
Rk51	net4#13	net4#14	0.903764	$metal1_conn
Rk52	net8#4	net8#5	37.511574	$metal1_conn
Rk53	net27	net27#2	0.168981	$metal1_conn
Rk55	net27#2	net27#5	0.745057	$metal1_conn
Rk56	net27#5	net27#7	0.002894	$metal1_conn
Rk57	net27#7	net27#8	0.157084	$metal1_conn
Rk58	net27#5	net27#9	0.152819	$metal1_conn
Rk59	net27#3	net27#2	15.500000	$metal1_conn
Rk60	net27#6	net27#7	15.500000	$metal1_conn
Rk61	net6#6	net6#7	75.000000	$metal1_conn
Rk62	net6#8	net6#9	31.001551	$metal1_conn
Rk63	PHI#5	PHI#8	47.069946	$metal1_conn
Rk64	PHI#8	PHI	0.231921	$metal1_conn
Rk65	net21	net21#2	37.504650	$metal1_conn
Rk66	net1#4	net1#5	0.158561	$metal1_conn
Rk67	net1#5	net1#7	0.005787	$metal1_conn
Rk68	net1#7	net1#8	0.167379	$metal1_conn
Rk69	net1#6	net1#7	15.500000	$metal1_conn
Rk70	net6#10	net6#11	0.916748	$metal1_conn
Rk71	VDD#21	VDD#22	0.149564	$metal1_conn
Rk72	VDD#22	VDD#24	0.011574	$metal1_conn
Rk73	VDD#24	VDD#25	0.166843	$metal1_conn
Rk74	VDD#23	VDD#24	15.500000	$metal1_conn
Rk75	net14	net14#2	0.160250	$metal1_conn
Rk76	net14#2	net14#4	0.002894	$metal1_conn
Rk77	net14#4	net14#5	0.164837	$metal1_conn
Rk78	net14#3	net14#4	15.500000	$metal1_conn
Rk79	GND#13	GND#14	37.501549	$metal1_conn
Rk80	GND#15	GND#16	75.002892	$metal1_conn
Rk81	net6#3	net6#13	45.424999	$metal1_conn
Rk82	net18	net18#2	0.153126	$metal1_conn
Rk83	net18#2	net18#4	0.008681	$metal1_conn
Rk84	net18#4	net18#5	0.166175	$metal1_conn
Rk85	net18#3	net18#4	15.500000	$metal1_conn
Rk86	net33#3	net33#4	37.504650	$metal1_conn
Rk87	COUT#1	COUT#2	75.002892	$metal1_conn
Rk88	COUT#3	COUT#4	0.160250	$metal1_conn
Rk89	COUT#4	COUT#6	0.002894	$metal1_conn
Rk90	COUT#6	COUT#7	0.164837	$metal1_conn
Rk91	COUT#5	COUT#6	15.500000	$metal1_conn
Rk92	net33#5	net33#6	1.199497	$metal1_conn
Rk93	GND#17	GND#18	75.002892	$metal1_conn
Rk94	VDD#26	VDD#27	31.001551	$metal1_conn
Rk95	VDD#28	VDD#29	0.163813	$metal1_conn
Rk97	VDD#29	VDD#32	0.164169	$metal1_conn
Rk98	VDD#30	VDD#29	15.500000	$metal1_conn
Rk99	GND#19	GND#20	37.501549	$metal1_conn
Rk100	SOUT#9	SOUT#10	75.002892	$metal1_conn
Rk101	SOUT#11	SOUT#12	31.251551	$metal1_conn
Rk102	net21#3	net21#4	37.503101	$metal1_conn
Rk103	net21#5	net21#6	1.195367	$metal1_conn
Rk104	SOUT#13	SOUT#14	0.324495	$metal1_conn
Rk105	SOUT#14	SOUT#15	2.577441	$metal1_conn
Rk106	GND#21	GND#22	75.000000	$metal1_conn
Rk107	VDD#33	VDD#34	0.153126	$metal1_conn
Rk108	VDD#34	VDD#36	0.008681	$metal1_conn
Rk109	VDD#36	VDD#37	0.166175	$metal1_conn
Rk110	VDD#35	VDD#36	15.500000	$metal1_conn
Rk111	SOUT#16	SOUT#17	0.103290	$metal1_conn
Rk112	SOUT#17	SOUT#5	46.499588	$metal1_conn
Rk113	net18#6	net18#7	0.160250	$metal1_conn
Rk114	net18#7	net18#9	0.002894	$metal1_conn
Rk115	net18#9	net18#10	0.164837	$metal1_conn
Rk116	net18#8	net18#9	15.500000	$metal1_conn
Rk117	net37#3	net37#4	37.501549	$metal1_conn
Rk118	net18#11	net18#12	0.615361	$metal1_conn
Rk119	net37#5	net37#6	2.409303	$metal1_conn
Rk120	net3#5	net3#12	46.248158	$metal1_conn
Rk121	net14#6	net14#8	0.164481	$metal1_conn
Rk122	net14#8	net14#9	0.002894	$metal1_conn
Rk123	net14#9	net14#10	0.160607	$metal1_conn
Rk124	net14#7	net14#8	15.500000	$metal1_conn
Rk125	COUT#8	COUT#9	75.000000	$metal1_conn
Rk126	net14#11	net14#12	0.859018	$metal1_conn
Rk127	net2#13	net2#14	0.146001	$metal1_conn
Rk128	net2#14	net2#16	0.014468	$metal1_conn
Rk129	net2#16	net2#17	0.167512	$metal1_conn
Rk130	net2#15	net2#16	15.500000	$metal1_conn
Rk131	net2#18	net2#19	2.400260	$metal1_conn
Rk132	net2#19	net2#20	1.220229	$metal1_conn
Rk133	net2#21	net2#22	37.501549	$metal1_conn
Rk134	net1#9	net1#10	1.663371	$metal1_conn
Rk135	net1#11	net1#2	46.186584	$metal1_conn
Rk136	net5	net5#2	0.149899	$metal1_conn
Rk137	net5#2	net5#4	0.006430	$metal1_conn
Rk138	net5#2	net5#6	0.811109	$metal1_conn
Rk140	net5#4	net5#8	0.156788	$metal1_conn
Rk141	net5#6	net5#9	0.149613	$metal1_conn
Rk142	net5#6	net5#10	0.157075	$metal1_conn
Rk143	net5#3	net5#4	15.500000	$metal1_conn
Rk144	net5#5	net5#6	15.500000	$metal1_conn
Rk145	net1#13	net1#15	0.187877	$metal1_conn
Rk147	net1#14	net1#15	37.500000	$metal1_conn
Rk148	CIN#5	CIN#8	45.436287	$metal1_conn
Rk149	CIN	CIN#9	0.463466	$metal1_conn
Rk150	CIN#9	CIN#10	3.391644	$metal1_conn
Rk151	net7#2	net7#9	49.371017	$metal1_conn
Rk152	net12#3	net12#4	37.503101	$metal1_conn
Rk153	net12#5	net12#6	2.908509	$metal1_conn
Rk154	net3#13	net3#14	3.842346	$metal1_conn
Rk155	net3#15	net3#16	2.083880	$metal1_conn
Rk156	net3#16	net3#2	45.548016	$metal1_conn
Rk157	COUT#10	COUT#11	0.704036	$metal1_conn
Rk158	COUT#11	COUT#12	1.228367	$metal1_conn
Rk159	net8#6	net8#2	46.737949	$metal1_conn
Rk160	net8#8	net8#9	0.149256	$metal1_conn
Rk161	net8#9	net8#11	0.006430	$metal1_conn
Rk162	net8#11	net8#12	0.157431	$metal1_conn
Rk163	net8#9	net8#13	1.080681	$metal1_conn
Rk164	net8#10	net8#11	15.500000	$metal1_conn
Rk165	net8#14	net8#15	2.680126	$metal1_conn
Rk166	VDD#38	VDD	0.299241	$metal1_conn
Rk167	VDD	VDD#39	0.122606	$metal1_conn
Rk168	VDD#39	VDD#40	0.167150	$metal1_conn
Rk169	VDD#40	VDD#42	0.172346	$metal1_conn
Rk170	VDD#42	VDD#43	0.198321	$metal1_conn
Rk171	VDD#43	VDD#44	0.207410	$metal1_conn
Rk172	VDD#44	VDD#45	0.072207	$metal1_conn
Rk173	VDD#45	VDD#46	0.240793	$metal1_conn
Rk174	VDD#41	VDD#42	18.750000	$metal1_conn
Rk175	GND#23	GND	0.242094	$metal1_conn
Rk176	GND	GND#24	0.387296	$metal1_conn
Rk177	GND#24	GND#26	0.377944	$metal1_conn
Rk178	GND#26	GND#27	0.200533	$metal1_conn
Rk179	GND#27	GND#28	0.313787	$metal1_conn
Rk180	GND#25	GND#26	15.500000	$metal1_conn
Rk181	VDD#47	VDD	0.389636	$metal1_conn
Rk182	VDD	VDD#49	0.128840	$metal1_conn
Rk183	VDD#49	VDD#50	0.076888	$metal1_conn
Rk184	VDD#50	VDD#51	0.064719	$metal1_conn
Rk185	VDD#51	VDD#52	0.266158	$metal1_conn
Rk186	VDD#52	VDD#53	0.312106	$metal1_conn
Rk187	VDD#53	VDD#54	0.030662	$metal1_conn
Rk188	VDD#48	VDD#49	18.750000	$metal1_conn
Rk189	GND#29	GND	0.863661	$metal1_conn
Rk190	GND	GND#30	0.099747	$metal1_conn
Rk191	GND#30	GND#32	0.116371	$metal1_conn
Rk192	GND#32	GND#33	0.120527	$metal1_conn
Rk193	GND#33	GND#34	0.300280	$metal1_conn
Rk194	GND#34	GND#35	0.278198	$metal1_conn
Rk195	GND#35	GND#36	0.354047	$metal1_conn
Rk196	GND#31	GND#32	15.500000	$metal1_conn
Rk197	GND#37	GND	0.286772	$metal1_conn
Rk198	GND	GND#38	0.348075	$metal1_conn
Rk199	GND#38	GND#40	0.167284	$metal1_conn
Rk200	GND#40	GND#41	0.165206	$metal1_conn
Rk201	GND#41	GND#42	0.343919	$metal1_conn
Rk202	GND#39	GND#40	15.500000	$metal1_conn
Rk203	COUT	COUT#13	0.898066	$metal1_conn
Rk209	PHI#2	PHI#8	45.000000	$metal1_conn
Rk215	CIN#2	CIN#9	45.000000	$metal1_conn
Rj1	VDD#46	VDD#1	1.035883	$metal2_conn
Rj2	GND#1	GND#28	1.272682	$metal2_conn
Rj3	net7#5	net7#9	0.599605	$metal2_conn
Rj4	net7#9	net7#6	0.461924	$metal2_conn
Rj5	SOUT#8	SOUT#15	2.020458	$metal2_conn
Rj6	net2#20	net2#5	2.278064	$metal2_conn
Rj7	GND#42	GND#4	1.067352	$metal2_conn
Rj8	VDD#3	VDD#54	1.195370	$metal2_conn
Rj9	net10#6	net10	0.924778	$metal2_conn
Rj10	VDD#6	VDD#45	1.263018	$metal2_conn
Rj11	VDD#53	VDD#8	1.391929	$metal2_conn
Rj12	GND#5	GND#35	1.146224	$metal2_conn
Rj13	net3#7	net3#14	0.400648	$metal2_conn
Rj14	net3#14	net3#9	0.729194	$metal2_conn
Rj15	net4#4	net4#14	0.668794	$metal2_conn
Rj16	net4#14	net4#7	0.400618	$metal2_conn
Rj17	net37#2	net37#6	0.921536	$metal2_conn
Rj18	GND#8	GND#27	1.284842	$metal2_conn
Rj19	VDD#44	VDD#13	1.299584	$metal2_conn
Rj20	net12#2	net12#6	0.955360	$metal2_conn
Rj21	net4#13	net4#9	2.258736	$metal2_conn
Rj22	net33#6	net33	0.911474	$metal2_conn
Rj23	GND#34	GND#9	1.042489	$metal2_conn
Rj24	VDD#17	VDD#43	1.267880	$metal2_conn
Rj25	GND#41	GND#11	1.057627	$metal2_conn
Rj26	VDD#20	VDD#52	1.185706	$metal2_conn
Rj27	net2#25	net2#7	0.614847	$metal2_conn
Rj28	net2#25	net2#9	0.705701	$metal2_conn
Rj29	net10#5	net10#3	0.926154	$metal2_conn
Rj30	net4#12	net4#11	0.900648	$metal2_conn
Rj31	net8#4	net8#15	1.099311	$metal2_conn
Rj32	net6#7	net6#11	0.620443	$metal2_conn
Rj33	net6#11	net6#9	0.511754	$metal2_conn
Rj34	net21	net21#6	1.021571	$metal2_conn
Rj35	net1#10	net1#5	1.190864	$metal2_conn
Rj36	net3#16	net3#12	2.462485	$metal2_conn
Rj37	net6#10	net6#13	3.387813	$metal2_conn
Rj38	VDD#51	VDD#22	1.380015	$metal2_conn
Rj39	GND#14	GND#56	0.642095	$metal2_conn
Rj40	GND#56	GND#16	0.632615	$metal2_conn
Rj41	net14#2	net14#12	1.229520	$metal2_conn
Rj42	net18#12	net18#2	1.220192	$metal2_conn
Rj43	net33#5	net33#3	0.943983	$metal2_conn
Rj44	COUT#1	COUT#12	0.391015	$metal2_conn
Rj45	COUT#12	COUT#4	0.888450	$metal2_conn
Rj46	GND#38	GND#17	1.057658	$metal2_conn
Rj47	VDD#26	VDD#50	1.196287	$metal2_conn
Rj48	VDD#40	VDD#29	1.312428	$metal2_conn
Rj49	GND#19	GND#24	1.242864	$metal2_conn
Rj50	SOUT#9	SOUT#11	0.882227	$metal2_conn
Rj51	SOUT#11	SOUT#14	0.800930	$metal2_conn
Rj52	net21#3	net21#5	1.008512	$metal2_conn
Rj53	SOUT	SOUT#24	1.012304	$metal2_conn
Rj54	SOUT#24	SOUT#13	0.946960	$metal2_conn
Rj55	GND#30	GND#22	1.091482	$metal2_conn
Rj56	VDD#34	VDD#39	1.530962	$metal2_conn
Rj57	net18#11	net18#7	1.223325	$metal2_conn
Rj58	net37#4	net37#5	0.919946	$metal2_conn
Rj59	COUT#9	COUT#11	0.876458	$metal2_conn
Rj60	net14#9	net14#11	1.225493	$metal2_conn
Rj61	net2#14	net2#18	0.712151	$metal2_conn
Rj62	net2#18	net2#22	0.616959	$metal2_conn
Rj63	net1#9	net1#11	0.908304	$metal2_conn
Rj64	net1#11	net1#13	0.855152	$metal2_conn
Rj65	CIN#10	CIN#8	2.689690	$metal2_conn
Rj66	net12#3	net12#5	0.945696	$metal2_conn
Rj67	net3#13	net3#15	2.443616	$metal2_conn
Rj68	COUT#10	COUT#13	3.532706	$metal2_conn
Rj69	net8#6	net8#13	4.520224	$metal2_conn
Rj70	net8#13	net8#14	1.389088	$metal2_conn
Rj71	VDD#38	VDD#47	3.963225	$metal2_conn
Rj72	GND#37	GND#29	3.450795	$metal2_conn
Rj73	GND#29	GND#23	3.409021	$metal2_conn
Rj175	SOUT#17	SOUT#24	0.500000	$metal2_conn
Rj150	GND#33	GND#56	0.500000	$metal2_conn
Rj126	net2#19	net2#25	0.500000	$metal2_conn
*
*       CAPACITOR CARDS
*
*
C1	net27#9	VDD#44	5.95458e-18
C2	net6#10	SOUT#14	1.85058e-17
C3	net18#2	net18#3	6.5943e-18
C4	net33#5	net2#18	1.20574e-18
C5	GND#8	GND#7	9.2133e-18
C6	COUT#4	net6#5	4.9547e-18
C7	net4#14	RST#2	6.81544e-18
C8	SOUT#13	SOUT#17	4.3021e-18
C9	net14#3	COUT#4	2.16641e-17
C10	net4#2	net27#8	1.08666e-17
C11	SOUT#16	net8#2	5.4736e-18
C12	net4#11	net4#12	1.06847e-17
C13	VDD#25	net18#5	7.23963e-18
C14	net12#5	net1#13	1.21091e-17
C15	SOUT#14	SOUT#6	2.88521e-18
C16	net37#2	net2#20	5.58763e-18
C17	net21#3	net21#4	7.86296e-18
C18	net1#13	net7#3	1.28693e-18
C19	net18#12	net6	3.89547e-19
C20	net5#8	net5#3	5.41954e-18
C21	VDD#29	net5#10	1.56962e-18
C22	net2#12	net2#10	2.42848e-18
C23	net14	net3#12	1.17708e-17
C24	VDD#3	VDD#4	6.90574e-18
C25	net14#9	VDD#37	4.75174e-19
C26	VDD#3	CIN#3	6.5361e-18
C27	GND#11	SOUT#4	7.83961e-18
C28	VDD#32	net5#9	6.67107e-18
C29	net14#12	net3#6	4.15801e-19
C30	GND#28	PHI#3	1.48373e-18
C31	net2#18	net3#15	6.97617e-17
C32	net27	net27#3	6.4597e-18
C33	SOUT#8	net13#6	3.99894e-19
C34	net12#5	net1#3	4.02484e-18
C35	net2#18	net18#12	6.08839e-18
C36	net13	net13#3	3.4113e-18
C37	GND#41	SOUT#4	2.30176e-18
C38	VDD#45	net4#7	1.20264e-18
C39	VDD#44	net4#2	9.46832e-19
C40	net4#7	net4#6	9.11187e-18
C41	net21	net1#8	1.2762e-18
C42	GND#1	PHI#3	6.37645e-18
C43	net3#5	COUT#12	1.86334e-17
C44	net3#13	net8	1.31876e-17
C45	net18#2	net18	2.74444e-18
C46	net10#3	RST#1	7.10774e-18
C47	net3#12	net6#13	3.83023e-17
C48	VDD#41	net14#12	2.59275e-18
C49	COUT#4	COUT#5	1.1635e-17
C50	net10#5	RST#1	1.78681e-18
C51	VDD#40	net14#11	1.36899e-18
C52	VDD#26	net8#3	6.58737e-18
C53	net6#13	net18#5	5.08666e-19
C54	net4#12	net10#3	5.38967e-18
C55	net2#20	VDD#11	1.11731e-17
C56	net1#5	net1#4	1.02489e-18
C57	VDD#6	net4#7	5.73546e-17
C58	net18#8	net2#17	6.34564e-19
C59	net7#6	PHI#3	6.83721e-18
C60	VDD#20	net6#9	5.73546e-17
C61	net3#16	net33#6	3.83218e-17
C62	net4#11	net4#10	4.36387e-18
C63	net6#13	net3#16	1.55454e-16
C64	GND#34	net33	4.10975e-18
C65	net13#9	net13#3	2.02912e-18
C66	net12#5	net7#3	3.95976e-18
C67	net5	net8#8	7.12591e-18
C68	VDD#48	SOUT#13	1.85444e-17
C69	VDD#45	net2#3	2.32554e-18
C70	net18#12	VDD#50	2.01888e-17
C71	net2#20	SOUT#1	2.75641e-17
C72	GND#22	GND#30	3.33556e-18
C73	net12#3	net7#3	6.91777e-18
C74	net2#2	RST#1	6.90286e-19
C75	net4#9	net4#2	3.59209e-18
C76	net18#12	VDD#48	9.97543e-18
C77	COUT#10	net3#4	1.9504e-18
C78	net7#5	net4	1.61e-18
C79	net7#2	net5#8	5.45092e-18
C80	COUT#4	COUT#3	3.14327e-18
C81	VDD#6	net2#3	6.66865e-18
C82	net7#2	net1#2	6.24282e-17
C83	net18#3	net18#8	2.0708e-18
C84	SOUT#14	net8#3	1.85546e-18
C85	SOUT#14	SOUT#5	9.28904e-18
C86	net2#22	net2#21	5.54062e-18
C87	VDD#53	net3#9	3.82873e-18
C88	net18	net18#12	9.60203e-18
C89	net21#5	net12#6	1.10866e-17
C90	net14#12	COUT#7	9.1277e-18
C91	COUT#10	CIN#6	1.43083e-18
C92	net14#12	net3#12	3.81369e-18
C93	SOUT#11	net8#3	7.06242e-18
C94	net3#9	CIN#3	7.84181e-18
C95	VDD#29	net1	1.74901e-18
C96	net33	net2#7	5.80278e-17
C97	GND#5	GND#6	7.34192e-18
C98	VDD#40	net1	2.92742e-18
C99	net2#18	net2#17	1.50328e-17
C100	net8#15	PHI#6	1.4509e-18
C101	VDD#34	net6#5	1.40653e-18
C102	PHI#5	net4#3	1.23236e-17
C103	net2#20	net13#6	1.41333e-17
C104	net8#4	net8#5	3.3072e-18
C105	CIN#8	net3#15	1.67666e-16
C106	net10#3	net10#5	7.94554e-18
C107	net1#10	net1#4	1.18398e-17
C108	net8#14	net7#3	3.41523e-18
C109	net8#4	PHI#6	6.03822e-18
C110	net2#19	net2#12	1.33046e-17
C111	GND#8	PHI#5	4.8732e-18
C112	net10#6	GND#34	8.14279e-18
C113	net6#7	SOUT#4	8.73964e-18
C114	SOUT#17	net8#3	1.09923e-17
C115	net1#11	net5#8	2.21573e-18
C116	net4#7	net4#13	8.57949e-18
C117	VDD#33	net14#6	5.9888e-18
C118	CIN#10	net3#15	6.41882e-18
C119	net2#7	net33#6	3.14465e-17
C120	VDD#51	SOUT#14	4.75012e-17
C121	net12#2	net7#9	1.27311e-18
C122	VDD#8	SOUT#1	3.80632e-18
C123	VDD#20	CIN#2	3.48733e-18
C124	net6#7	net3#14	2.40277e-17
C125	VDD#30	PHI#4	1.18606e-18
C126	VDD#33	net3#5	1.11523e-17
C127	net12#5	net12#3	4.17429e-18
C128	CIN#10	net3#13	2.69246e-16
C129	net2#13	net2#15	5.37287e-18
C130	VDD#53	SOUT#1	2.357e-18
C131	net3#12	GND#16	1.36623e-17
C132	net3#12	RST#1	2.53357e-18
C133	net33#6	net3#2	3.44769e-17
C134	net2#8	VDD#52	2.46394e-18
C135	GND#11	net6#7	6.13228e-17
C136	net18#2	net18#8	1.05046e-18
C137	net6#13	VDD#23	2.08433e-18
C138	net14#2	COUT#7	8.96923e-19
C139	net14#3	net6#5	4.44372e-18
C140	GND#25	net8#15	4.06774e-17
C141	net4#7	net2#3	4.77177e-18
C142	net4#13	RST#2	4.26734e-17
C143	GND#30	net37#5	1.98627e-17
C144	net4#14	net4#13	4.81454e-18
C145	net2#7	net2#6	1.03847e-17
C146	CIN#10	COUT#13	4.94891e-18
C147	net33#6	net2#19	6.98998e-18
C148	net4#14	net2#3	6.6601e-18
C149	net1#11	net5#9	1.11583e-18
C150	CIN#8	COUT#10	6.12354e-18
C151	GND#28	net7#6	3.81828e-18
C152	GND#16	GND#15	5.52802e-18
C153	net18	net18#6	4.81107e-19
C154	net3#12	GND#34	1.14427e-17
C155	SOUT#11	net8#2	9.7462e-18
C156	net10	net4#4	5.72462e-17
C157	net12#6	PHI#5	2.6878e-17
C158	net4#9	net27	1.45032e-18
C159	VDD#26	VDD#27	8.5607e-18
C160	net3#12	GND#33	4.441e-18
C161	net1#9	net5	1.89372e-18
C162	net6#7	GND#41	7.97687e-18
C163	net12#2	PHI#5	1.42452e-17
C164	net2#17	net2#15	2.49227e-18
C165	GND#8	net12#6	2.65231e-17
C166	VDD#34	net3#6	3.78758e-18
C167	GND#4	CIN#1	7.83157e-18
C168	net2#18	net6	2.02439e-17
C169	net27#9	net4	1.60343e-18
C170	net13	SOUT#1	5.32049e-19
C171	net3#16	GND#34	4.61043e-18
C172	net6#13	GND#16	2.19708e-18
C173	net18#2	VDD#21	6.47808e-19
C174	net3#16	GND#33	3.58056e-18
C175	VDD#23	net6	3.74024e-18
C176	net5#8	net8#12	7.9977e-18
C177	net4#4	net10#6	1.084e-17
C178	net27#8	net4	1.66237e-18
C179	GND#1	net7#6	5.74685e-17
C180	net13#9	SOUT#1	5.98355e-19
C181	GND#1	PHI#2	2.08019e-17
C182	net14#6	net14#7	3.1048e-18
C183	GND#42	CIN#1	2.81595e-18
C184	GND#16	RST#1	1.22185e-18
C185	net4#9	net27#9	1.38655e-18
C186	PHI#5	net1#3	1.15731e-18
C187	net4#9	PHI#5	1.72164e-18
C188	net5#10	net1#9	1.22748e-17
C189	GND#19	net7#2	8.41408e-18
C190	net13#8	SOUT#1	1.05318e-18
C191	net7#9	net4#9	2.0581e-17
C192	net18#3	net6	3.24889e-18
C193	net8#8	VDD	5.38283e-18
C194	net14#11	net3#6	4.72163e-18
C195	net7#6	net4#3	1.70037e-18
C196	VDD#34	net14#6	6.82268e-19
C197	VDD#17	RST#2	1.37638e-18
C198	PHI#2	VDD#1	3.18312e-18
C199	GND#27	net12#6	1.15846e-17
C200	GND#8	net12#2	5.88321e-17
C201	net2	RST#1	4.37651e-19
C202	net14#9	net3#6	6.02364e-19
C203	net2#7	net3#16	6.52402e-18
C204	net3#15	COUT#13	4.61597e-17
C205	net8#14	net12#5	6.50915e-17
C206	net18#7	CIN#4	3.79893e-19
C207	net6#13	GND#33	6.22748e-17
C208	net6#2	CIN#5	1.95213e-18
C209	net3#12	net6#4	2.18531e-18
C210	CIN#10	net8#6	4.26282e-17
C211	net5	VDD	5.38283e-18
C212	RST#2	GND#9	5.69138e-18
C213	net18#11	CIN#4	6.01056e-19
C214	net2#18	net18#10	1.21911e-17
C215	CIN#8	net2#15	2.22697e-18
C216	net21#3	net1#2	9.06753e-19
C217	net2#19	net3#2	6.31571e-17
C218	net37#5	net37#4	1.02763e-17
C219	SOUT#17	net8#2	7.17818e-17
C220	net6#13	VDD#25	1.96834e-18
C221	VDD#34	net14#10	6.97776e-19
C222	net4#9	net27#8	2.2663e-18
C223	net2#13	VDD	4.03217e-18
C224	GND#17	GND#38	4.11518e-18
C225	net3#13	COUT#13	7.51707e-17
C226	GND#30	net6#3	3.25202e-18
C227	net3#15	COUT#10	2.42088e-17
C228	net12#3	net8#14	6.14727e-18
C229	net2#5	net10	1.70846e-17
C230	net14#6	VDD	3.88163e-18
C231	net7#6	PHI#2	2.44739e-17
C232	net14#10	net14#7	2.52549e-18
C233	SOUT#15	VDD#8	3.65712e-18
C234	COUT#4	net14	1.33445e-18
C235	net1#9	net1	5.20774e-18
C236	VDD#40	net1#9	5.55017e-17
C237	net3#16	net2#19	9.8947e-17
C238	net6#13	GND#14	1.35114e-17
C239	VDD#37	net14#10	6.02833e-18
C240	net14#2	net14#3	4.95248e-18
C241	SOUT#16	VDD	7.03798e-18
C242	net18#8	net6	8.15715e-19
C243	net8#4	net7#9	1.3668e-18
C244	VDD#34	VDD#35	9.00896e-18
C245	net3#16	net37#5	1.13856e-17
C246	VDD#39	net14#11	1.56252e-17
C247	net37#6	net33	8.91409e-18
C248	COUT#11	GND#22	2.47095e-17
C249	net18#7	net18#3	9.52773e-19
C250	net3#16	net6#2	1.40016e-18
C251	net2#18	CIN#4	1.54343e-17
C252	VDD#52	SOUT#14	6.43129e-17
C253	COUT#3	COUT#5	3.72954e-18
C254	net27	net1#8	7.69447e-18
C255	net7#9	PHI#2	1.68776e-16
C256	net2#8	net3	1.61265e-18
C257	net3#13	GND#39	4.07521e-18
C258	net6#13	net6#2	2.70865e-18
C259	net10	net2	6.48362e-18
C260	VDD#17	VDD#18	8.74142e-18
C261	net14#12	net14#5	1.03897e-17
C262	net14	VDD	3.74778e-18
C263	net12#2	net12	3.39271e-18
C264	GND#4	GND#42	4.05951e-18
C265	net6#13	net37#5	1.02187e-17
C266	VDD#34	net14#11	4.67193e-17
C267	net2#19	net13#9	1.18348e-17
C268	GND#31	net37#5	2.34961e-17
C269	net6#13	VDD#22	3.14196e-18
C270	net2#12	net3	1.67859e-18
C271	COUT#11	GND#30	4.58606e-18
C272	net2#5	net10#6	1.28092e-17
C273	net6#13	net2#19	2.35603e-17
C274	VDD#13	net4	1.53572e-18
C275	GND#22	COUT#9	5.7463e-17
C276	SOUT#8	VDD#8	7.86519e-18
C277	VDD#1	net7#5	6.39295e-17
C278	COUT#12	net3#12	2.59761e-17
C279	net6#7	net6#6	2.72909e-18
C280	GND#16	net6#4	8.41409e-18
C281	net10#6	net2	1.59515e-18
C282	net21	net1#3	2.11513e-18
C283	VDD#53	SOUT#15	6.16732e-17
C284	net2#7	GND#34	1.63187e-18
C285	VDD#12	net4	1.59419e-18
C286	net1#8	VDD	4.31456e-18
C287	net18#5	net18#10	5.46123e-19
C288	VDD#44	net4	3.95281e-18
C289	GND#14	GND#13	1.09819e-17
C290	SOUT#14	VDD#20	3.80992e-18
C291	VDD#16	net4	1.69788e-18
C292	net1#11	net7	3.29019e-18
C293	net14	COUT#3	5.92261e-18
C294	net37#6	net33#6	9.58373e-18
C295	net4#7	RST#3	9.31194e-19
C296	net4#13	net4#11	1.39919e-18
C297	VDD#34	net14#9	3.01681e-17
C298	VDD#34	net14#7	2.56991e-17
C299	net21#3	net7#2	7.49402e-18
C300	COUT#9	GND#30	6.44381e-18
C301	net6#11	CIN#2	3.69869e-17
C302	net13	VDD#52	3.95741e-18
C303	net3#13	net8#6	2.03853e-17
C304	VDD#30	net5#10	1.26916e-18
C305	net3#14	net3#7	1.06847e-17
C306	net6#10	VDD#22	7.79479e-18
C307	net18#6	net18#8	3.67439e-18
C308	net4#4	GND#35	1.92613e-18
C309	net13	VDD	2.99823e-18
C310	VDD#30	net1	4.19171e-18
C311	net7#2	VDD#32	5.11944e-18
C312	VDD#7	net13#6	1.07256e-17
C313	net13#9	VDD	3.50686e-18
C314	net8#15	net12#6	1.78933e-17
C315	net3#14	CIN#1	1.87042e-18
C316	net21#3	net1#13	7.62435e-18
C317	VDD#50	SOUT#14	4.73371e-17
C318	net13#8	VDD	2.8562e-18
C319	COUT#7	COUT#5	5.23184e-18
C320	net4#9	net4	1.29901e-18
C321	COUT#10	net8#13	5.38464e-17
C322	COUT#13	net8#6	1.69776e-16
C323	GND#33	net6#2	1.45199e-18
C324	net3#7	CIN#1	7.84713e-18
C325	net7#5	VDD#46	8.20379e-18
C326	VDD#20	SOUT#5	7.26379e-18
C327	VDD#14	net27#9	9.16617e-19
C328	GND#14	net6#2	8.26391e-18
C329	net4#13	net4#12	2.36682e-18
C330	COUT#12	net6#4	5.75204e-18
C331	net2#19	net13#6	7.58305e-18
C332	net6#10	VDD#51	4.0158e-17
C333	COUT#10	net8#6	5.60501e-17
C334	SOUT#14	VDD#26	1.67328e-17
C335	net14#2	net14#5	1.79038e-18
C336	COUT#1	net6#4	5.59846e-18
C337	VDD#52	net6#10	7.72908e-18
C338	GND#30	net2#22	3.49278e-18
C339	GND#35	net37#6	2.09743e-17
C340	net8#4	net12#6	1.16762e-17
C341	GND#19	GND#20	4.25438e-18
C342	net18#10	net18#8	5.43185e-18
C343	COUT#13	VDD#47	2.6128e-17
C344	net18#7	net2#13	9.13245e-19
C345	GND#19	net12#5	1.48301e-17
C346	GND#24	net8#15	9.54758e-17
C347	net12#6	net12#2	7.2986e-18
C348	VDD#41	VDD	5.04836e-17
C349	VDD#13	net4#9	5.24004e-18
C350	net4#12	RST#2	2.79498e-17
C351	VDD#11	net13#6	3.92427e-18
C352	VDD#26	SOUT#11	7.22437e-17
C353	COUT#3	net6#5	1.37307e-18
C354	net18#10	net6	4.85417e-19
C355	GND#5	SOUT#3	6.89827e-18
C356	GND#8	PHI#3	1.66757e-18
C357	net8#13	net7	1.69935e-18
C358	VDD#20	net6#10	7.18163e-18
C359	COUT#7	net6#5	1.51638e-18
C360	VDD#48	VDD	1.84109e-17
C361	VDD#14	net27#8	8.71787e-19
C362	PHI#4	net1#2	8.74316e-19
C363	net3#13	GND#17	1.34681e-17
C364	net33#3	net6#2	5.33847e-18
C365	net12#6	net7#2	1.17173e-17
C366	net8#15	net21#6	1.08881e-16
C367	net8#13	VDD#38	2.41494e-16
C368	GND#33	net37#5	2.14797e-17
C369	COUT#1	GND#22	1.03409e-17
C370	GND#5	net37#6	1.81945e-17
C371	net1#4	PHI#4	1.44489e-18
C372	RST#2	net10#5	9.80704e-18
C373	net33#5	net6#2	1.07286e-17
C374	net14#11	net3#5	9.08769e-18
C375	net27#9	net27#6	4.75038e-18
C376	net18#3	CIN#4	8.11298e-19
C377	net14#7	net3#6	3.21061e-18
C378	net6#13	net33#3	2.51269e-18
C379	net1#8	PHI#4	1.88143e-18
C380	net4#9	VDD#44	2.06922e-17
C381	net3#13	GND#38	1.313e-17
C382	net3#16	net33#5	7.58749e-17
C383	net4#4	net2	5.30553e-18
C384	SOUT#9	CIN#10	8.38618e-18
C385	net4#13	RST#3	7.58286e-19
C386	net13#6	VDD	2.25483e-17
C387	net2#5	net2#2	2.35794e-18
C388	net8#13	VDD#47	2.50154e-17
C389	VDD#3	CIN#2	4.70316e-18
C390	GND#23	net8#14	5.33993e-17
C391	COUT#10	GND#29	1.71437e-17
C392	COUT#13	GND#37	3.86048e-18
C393	net2#5	GND#35	5.74691e-17
C394	GND#14	net37#5	2.82455e-17
C395	net18#6	net2#13	5.19581e-18
C396	net3#14	GND#39	1.07545e-17
C397	net6#9	net6#8	8.08013e-18
C398	net18#7	net18#8	9.88123e-18
C399	SOUT#15	net3#9	5.92466e-18
C400	net14	net6#5	1.61265e-18
C401	GND#17	SOUT#9	5.73546e-17
C402	net3#5	COUT#11	1.75417e-17
C403	net8#8	net8#10	6.1458e-18
C404	CIN#2	GND#4	7.43834e-18
C405	net8#6	VDD#47	2.00796e-16
C406	net8#13	GND#23	5.72913e-17
C407	net14#5	net6#5	1.67859e-18
C408	net14#3	VDD	1.63389e-18
C409	VDD#8	VDD#9	1.00973e-17
C410	net6#13	net33#5	1.57779e-17
C411	net18#7	net2#14	1.99961e-17
C412	GND#5	net37#2	5.94147e-17
C413	net18#11	net2#13	5.69125e-19
C414	net37#4	net2#22	5.90816e-17
C415	net14#5	COUT#7	6.35918e-18
C416	net2#9	net6#13	5.82886e-18
C417	VDD#43	net4#11	3.22088e-18
C418	VDD#43	RST#3	1.47631e-18
C419	GND#19	PHI#6	2.13222e-18
C420	net2#19	net3	7.70154e-18
C421	net27	PHI#4	1.65648e-18
C422	net18#8	CIN#4	2.90806e-18
C423	net21#6	GND#25	1.93046e-18
C424	net5#10	net1	1.88143e-18
C425	net8#13	GND#29	2.34639e-17
C426	VDD#17	RST#3	5.84522e-18
C427	net6#10	CIN#2	2.2978e-17
C428	net7#9	VDD#16	4.7682e-18
C429	SOUT#9	GND#38	7.98287e-18
C430	net14#7	VDD	1.76681e-18
C431	net6#10	net3#14	1.82188e-18
C432	net5#9	net1	1.6651e-18
C433	net27#8	net27#6	4.25234e-18
C434	net7#9	net4#2	3.86949e-17
C435	net12#3	net8#10	1.36416e-18
C436	net2#15	CIN#4	3.36679e-18
C437	net14#9	COUT#11	1.85386e-18
C438	net8#4	net21	6.53006e-17
C439	net18#6	net2#15	6.34565e-19
C440	net2#20	GND#35	5.51468e-18
C441	net37#4	net2#18	9.96159e-19
C442	VDD#1	VDD	2.00865e-17
C443	net5#10	net5#5	5.98337e-18
C444	GND#23	VDD#38	1.68965e-17
C445	VDD#46	VDD	9.5977e-17
C446	net10#3	net3#12	8.30508e-18
C447	net18	net6	1.29063e-18
C448	net7#5	VDD	1.83234e-17
C449	net21	net21#2	5.56319e-18
C450	net6#13	net18#2	7.94215e-19
C451	net18#7	net2#15	1.51212e-18
C452	net7#9	VDD	8.68679e-18
C453	net1#9	VDD#39	6.60386e-17
C454	SOUT#2	net2#20	1.99233e-17
C455	SOUT#15	VDD	1.1934e-16
C456	SOUT#8	VDD	2.60209e-17
C457	net18#5	net6	1.57665e-18
C458	VDD#17	net4#11	6.26705e-17
C459	net2#9	net6#10	2.25842e-18
C460	VDD#22	net18	6.19933e-19
C461	COUT#4	net3#12	1.46298e-17
C462	SOUT#5	CIN#10	1.30767e-17
C463	net8#12	net8#10	5.02791e-18
C464	net4#7	net4#14	7.36443e-18
C465	net2#20	VDD	4.57679e-17
C466	net37#4	net37#3	5.72918e-18
C467	net4#9	PHI#4	6.03374e-18
C468	VDD#54	VDD	1.23253e-16
C469	VDD#3	VDD	2.7857e-17
C470	VDD#38	GND#29	2.92267e-16
C471	net8#6	GND#37	5.14604e-17
C472	net14	net14#3	6.43098e-18
C473	VDD#22	VDD#23	6.83853e-18
C474	net2#9	net3	5.04571e-18
C475	net18#7	net2#18	4.44358e-19
C476	VDD#45	VDD	7.75233e-17
C477	net1#11	net1#2	1.30301e-18
C478	SOUT#13	CIN#10	1.01282e-17
C479	VDD#6	VDD	2.73683e-17
C480	net18#8	net2#15	2.42745e-17
C481	net2#22	CIN#5	2.01578e-17
C482	GND#17	net8	7.41976e-18
C483	net6#9	SOUT#5	1.42367e-17
C484	GND#16	COUT#1	6.53236e-17
C485	net18	net18#3	3.40485e-18
C486	VDD#53	VDD	4.18757e-17
C487	net8#4	PHI#5	1.36376e-17
C488	net10#5	net3#12	4.39577e-18
C489	VDD#47	GND#29	2.87781e-16
C490	net21#5	net12#5	1.10373e-16
C491	net1#2	net1#9	2.72292e-18
C492	net3#9	VDD	1.57428e-17
C493	net18#2	net18#6	5.26452e-19
C494	COUT#11	COUT#9	1.24425e-17
C495	GND#34	net37#6	4.55157e-17
C496	net2#18	net18#11	7.86867e-18
C497	net2#20	GND#5	3.03104e-17
C498	net4#7	VDD	7.05558e-18
C499	net6#11	SOUT#5	4.10628e-17
C500	GND#24	net8#14	2.12408e-17
C501	SOUT#17	CIN#10	3.89817e-17
C502	net4#14	VDD	1.9938e-17
C503	VDD#17	net4#12	1.3639e-17
C504	net5#9	net5#5	5.24259e-18
C505	net37#5	net33#6	8.7882e-19
C506	GND#37	VDD#47	2.4242e-17
C507	VDD#21	net6	1.49699e-18
C508	VDD#23	net18#3	2.67659e-17
C509	net12#5	net21#3	7.27979e-18
C510	VDD#13	VDD	8.59973e-18
C511	net2#18	net18#5	1.11731e-17
C512	COUT#1	GND#33	6.41545e-18
C513	VDD#44	VDD	5.01915e-17
C514	VDD#25	net6	1.76343e-18
C515	net7#2	net1#8	3.56475e-18
C516	net18#7	net18#6	1.52878e-18
C517	net12#3	net8#12	3.48692e-18
C518	net4#11	RST#3	7.27484e-18
C519	net2#20	net13#8	1.14928e-17
C520	net3#16	net37#6	2.48702e-18
C521	PHI#2	VDD#2	2.42465e-18
C522	net3#14	GND#11	1.13087e-17
C523	net6#10	net18#12	1.97795e-18
C524	net4#9	VDD	2.30143e-17
C525	net21	net7#9	2.53114e-18
C526	GND#24	net21#5	9.83093e-18
C527	net4#13	VDD	5.55753e-17
C528	VDD#20	SOUT#6	6.64336e-18
C529	net14#5	net14#3	3.55686e-18
C530	net2#3	RST#3	6.91892e-19
C531	net4#12	RST#3	1.09625e-17
C532	CIN#10	net8#2	1.29162e-16
C533	net2#2	net10	1.34514e-17
C534	net37#5	net33#3	1.28305e-17
C535	net1#13	net7#2	7.04502e-18
C536	SOUT#9	net3#13	1.96049e-17
C537	VDD#43	VDD	6.6263e-17
C538	VDD#26	SOUT#17	1.34037e-17
C539	GND#8	net4#3	6.92722e-18
C540	net2#19	VDD#25	1.11731e-17
C541	VDD#17	VDD	1.87066e-17
C542	net18#5	net18#3	5.62966e-18
C543	VDD#22	net18#3	1.36665e-18
C544	net37#6	net2#7	1.12161e-17
C545	net37#6	net3#3	3.45245e-18
C546	net3#2	net3#16	3.17639e-18
C547	net18#11	VDD#48	1.82285e-17
C548	net2#19	VDD	9.44797e-17
C549	VDD#52	VDD	7.34476e-17
C550	net1#11	net7#2	5.32192e-17
C551	VDD#45	net4#9	2.27516e-18
C552	GND#27	net4#3	2.34451e-18
C553	VDD#20	VDD	2.54215e-17
C554	net33#3	GND#33	1.43923e-18
C555	net2#2	net10#6	2.95457e-18
C556	net21#6	net12#6	1.20325e-16
C557	SOUT#14	SOUT#11	3.9452e-18
C558	COUT#1	COUT#2	2.43886e-18
C559	net37#2	net3#3	1.93734e-18
C560	GND#19	net21#5	1.60436e-17
C561	net4#11	VDD	1.33211e-17
C562	net37#5	net33#5	1.1788e-17
C563	net4#12	VDD	2.20512e-17
C564	net3#12	RST#2	9.91286e-18
C565	net13	net2#8	6.36784e-18
C566	VDD#8	net13#6	4.28628e-17
C567	net33#3	net37#4	1.03108e-17
C568	RST	net2#5	2.37099e-17
C569	net14#6	net3#6	1.6651e-18
C570	net18#10	net2#17	6.35916e-18
C571	net13	net2#9	1.06131e-18
C572	net3#14	SOUT#4	1.6268e-17
C573	net6#9	VDD	7.37058e-18
C574	net3#14	GND#41	1.66716e-17
C575	VDD#28	net1	1.62659e-18
C576	net3#16	net2#18	4.94495e-17
C577	SOUT#9	net8	7.97071e-18
C578	COUT#11	GND#31	2.26769e-18
C579	net4#4	RST#1	2.05029e-18
C580	net14#10	net3#6	1.61378e-18
C581	VDD#6	RST	5.82138e-18
C582	net10	RST	1.06575e-18
C583	VDD#32	net1	1.6651e-18
C584	RST	net10#6	2.54666e-18
C585	net1#5	VDD	7.26628e-18
C586	SOUT#14	net6#9	6.25922e-18
C587	GND#14	net33#3	5.84121e-17
C588	net1#10	VDD	5.70763e-17
C589	net3#12	VDD	6.00819e-17
C590	GND#19	net21#3	7.02068e-17
C591	GND#9	net10#3	6.14823e-17
C592	net3#16	VDD	1.44134e-17
C593	net6#13	VDD	6.92227e-18
C594	net3#9	CIN#2	4.08481e-18
C595	net6#10	VDD	3.28553e-17
C596	COUT#4	net14#12	6.63795e-19
C597	VDD#28	net1#9	1.04369e-17
C598	net14#12	VDD	3.97681e-17
C599	net4#14	RST	3.30628e-17
C600	net14#9	net14#7	5.30663e-18
C601	net6#10	VDD#50	5.9841e-18
C602	RST	net4#4	4.07578e-18
C603	net14#2	VDD	6.72049e-18
C604	net12#6	net21	7.43001e-18
C605	VDD#45	net4#13	8.3269e-18
C606	net18#11	net18#6	1.0426e-17
C607	VDD#51	VDD	5.07658e-17
C608	COUT#4	VDD#34	5.58455e-18
C609	net3#14	CIN#2	1.74974e-16
C610	net13#9	net2#9	1.88405e-18
C611	net14#11	net14#10	1.11682e-17
C612	SOUT#11	SOUT#12	8.05404e-18
C613	net8#8	net7	1.74376e-18
C614	VDD#48	SOUT#14	2.30344e-17
C615	GND#14	net33#5	9.51969e-18
C616	net18#12	VDD	2.30345e-17
C617	COUT#4	VDD	3.08743e-18
C618	net8#12	net7	1.89454e-18
C619	net2#9	VDD#52	3.31251e-18
C620	net6#9	SOUT#6	6.36586e-18
C621	VDD#50	VDD	1.60024e-17
C622	net14#2	COUT#4	2.04995e-17
C623	VDD#26	VDD	1.20899e-17
C624	net13#6	VDD#53	1.49759e-17
C625	net21#5	net1#3	9.17556e-19
C626	net1#10	VDD#41	8.85271e-17
C627	GND#9	net10#5	2.40058e-17
C628	net18#7	CIN#8	2.60427e-18
C629	net6#10	VDD#26	1.20141e-17
C630	VDD#29	VDD	9.1833e-18
C631	VDD#40	VDD	2.99529e-17
C632	net21#3	net1#3	7.56451e-18
C633	net10	net10#6	5.26313e-18
C634	SOUT#14	VDD	6.6719e-17
C635	GND#9	net2	1.84566e-18
C636	SOUT#17	net3#13	1.56232e-17
C637	net2#17	CIN#4	1.79524e-18
C638	SOUT#11	VDD	8.61553e-18
C639	net10	net10#2	7.36722e-18
C640	net13#6	SOUT#1	7.27353e-18
C641	VDD#6	net4#13	8.24438e-18
C642	VDD#3	net3#9	5.7463e-17
C643	net6#10	SOUT#5	4.85612e-17
C644	COUT#12	COUT#1	1.30153e-17
C645	net8#15	net21#5	8.01512e-17
C646	net12#5	net7#2	2.08289e-17
C647	SOUT#13	VDD	3.07007e-17
C648	net7#9	PHI#5	1.57736e-16
C649	net18#2	net18#7	2.47864e-18
C650	net18#11	CIN#8	7.28111e-18
C651	SOUT#17	VDD	3.95099e-17
C652	net33#3	net33#4	7.44269e-18
C653	net8#15	net12#5	1.51553e-17
C654	GND#17	SOUT	4.81382e-18
C655	net3#15	CIN#5	4.47454e-17
C656	VDD#39	VDD	4.81274e-17
C657	SOUT	GND#38	4.51982e-17
C658	net1#4	net1#6	3.58452e-18
C659	GND#11	GND#41	4.11518e-18
C660	net37#5	net6#2	1.56376e-17
C661	net18#7	VDD	7.8066e-19
C662	GND#34	net10#5	9.26507e-17
C663	net18#11	VDD	3.78618e-17
C664	COUT#3	net3#12	1.11869e-17
C665	GND#5	SOUT#2	1.00582e-17
C666	net14#11	VDD	3.508e-17
C667	SOUT#9	SOUT	3.26552e-18
C668	net14#9	VDD	6.51924e-18
C669	net37#4	net6#2	1.17656e-18
C670	net5	net7	1.74376e-18
C671	net18#6	CIN#4	1.36381e-18
C672	net2#18	VDD	3.68935e-17
C673	VDD#22	net18#2	2.4189e-17
C674	SOUT#9	SOUT#10	4.02702e-18
C675	net5#8	net7	1.89454e-18
C676	net1#11	VDD	2.21495e-17
C677	net18#10	CIN#4	1.51804e-18
C678	net1#9	VDD	4.34033e-17
C679	VDD#37	net14#7	6.34561e-19
C680	net7#9	net27	4.7682e-18
C681	CIN#8	VDD	3.09461e-17
C682	net14#9	net14#10	1.54087e-18
C683	CIN#10	VDD	4.01705e-17
C684	GND#22	net3#4	5.30034e-18
C685	net33	net3#3	5.56036e-18
C686	SOUT#14	SOUT#13	8.24937e-18
C687	net1#5	PHI#4	4.59686e-18
C688	net3#15	VDD	6.9179e-17
C689	net3#13	VDD	2.12072e-17
C690	GND#8	PHI#2	9.37699e-18
C691	net18#12	net18#11	3.62642e-18
C692	COUT#13	VDD	4.05294e-17
C693	net4#14	net2#2	1.00706e-18
C694	net3#9	net3#10	7.78712e-18
C695	COUT#10	VDD	8.28361e-18
C696	VDD#14	net4	4.31944e-18
C697	net13#9	net2#12	6.35934e-18
C698	net33#6	net3#3	9.74256e-18
C699	net21	net1#6	9.87673e-19
C700	net13#6	net13	5.9474e-19
C701	net8#13	VDD	1.05209e-16
C702	net8#6	VDD	4.75508e-17
C703	VDD#22	net18#12	1.33526e-17
C704	net37#5	net3#15	6.87187e-18
C705	net1#8	net1#6	2.49885e-18
C706	VDD#38	VDD	1.08654e-16
C707	VDD#12	net27#9	5.92276e-18
C708	VDD#47	VDD	1.30247e-16
C709	net21#3	net7#3	1.24534e-18
C710	GND#23	VDD	4.10123e-17
C711	net1#10	VDD#40	2.64148e-17
C712	GND#29	VDD	1.03701e-16
C713	net12#3	net12#4	8.58427e-18
C714	GND#37	VDD	4.57179e-17
C715	net4#4	net2#2	5.9339e-18
C716	SOUT#11	SOUT#13	5.12065e-18
C717	PHI#2	VDD	9.91243e-18
C718	SOUT#14	SOUT#17	1.04139e-17
C719	CIN#2	VDD	9.27084e-18
C720	net2#14	net18#8	1.46766e-18
C721	SOUT#2	VDD	3.19199e-18
C722	GND#30	CIN#6	2.27489e-18
C723	net4#2	VDD	3.36886e-17
C724	net37#4	net3#15	6.69749e-18
C725	net3#2	VDD	1.39872e-17
C726	RST#2	VDD	4.89099e-18
C727	SOUT#2	net3#2	2.96414e-18
C728	VDD#21	net18	5.39378e-18
C729	net2#2	RST#2	4.68438e-19
C730	SOUT#5	VDD	4.71181e-17
C731	CIN#2	SOUT#5	2.24903e-17
C732	net37#6	net37#2	5.42102e-18
C733	PHI#5	VDD	3.92957e-18
C734	RST#2	net10#6	4.97058e-18
C735	net6#9	net6#10	1.28612e-17
C736	VDD#51	net18#12	1.58936e-17
C737	net1#2	VDD	4.05185e-17
C738	net8#13	net7#2	5.03908e-18
C739	VDD#41	PHI#4	4.00553e-18
C740	net3#5	VDD	5.23543e-17
C741	net3#12	net6#5	3.06697e-17
C742	CIN#5	VDD	3.59722e-18
C743	net14#6	COUT#11	4.02949e-18
C744	net7#2	VDD	1.55004e-17
C745	SOUT#11	SOUT#17	3.35024e-17
C746	net2#5	net4#4	8.60035e-18
C747	VDD#28	net5#10	6.09903e-18
C748	net2#14	CIN#8	6.74273e-18
C749	GND#16	net6#3	6.81271e-18
C750	net12#6	PHI#6	3.97093e-18
C751	RST	net2#2	3.581e-17
C752	VDD#52	SOUT#15	3.31388e-17
C753	net1#5	net1#6	3.82133e-18
C754	VDD#1	PHI#1	7.09794e-18
C755	net13#6	net13#9	4.5631e-19
C756	net10#3	net10#4	1.02675e-17
C757	net33	net33#6	6.38516e-18
C758	net12#2	PHI#6	1.88117e-18
C759	net33#3	net33#5	8.08775e-18
C760	net4#9	VDD#43	1.98786e-17
C761	VDD#46	PHI#1	2.34624e-18
C762	GND#33	net6#3	8.33848e-17
C763	GND#25	net12#6	2.42087e-17
C764	net1#2	net5#9	1.07149e-17
C765	net6#11	net6#10	7.96704e-18
C766	net18#5	CIN#4	5.0041e-19
C767	net2#14	net2#15	8.17507e-18
C768	SOUT#9	SOUT#17	1.72587e-17
C769	net14#12	net6#5	3.48736e-18
C770	net2#22	CIN#8	5.50796e-18
C771	net3#14	GND#42	1.10941e-17
C772	net2#7	net3#3	7.32354e-18
C773	PHI#1	VDD	3.08817e-17
C774	GND#4	net3#7	6.2996e-17
C775	CIN#3	VDD	2.28282e-17
C776	net14#2	net6#5	1.14794e-18
C777	net2#3	VDD	2.29897e-17
C778	SOUT#1	VDD	1.8004e-17
C779	net3#16	net6	1.04492e-17
C780	net4	VDD	1.0061e-17
C781	VDD#13	net27#9	1.39515e-18
C782	net7#5	PHI#1	8.89406e-18
C783	net3	VDD	1.18491e-17
C784	RST#3	VDD	1.72631e-17
C785	SOUT#6	VDD	1.04163e-17
C786	net21	net7#2	5.88649e-18
C787	GND#9	RST#1	5.7094e-18
C788	PHI#4	VDD	1.70111e-17
C789	COUT#11	net3#4	1.91864e-17
C790	net2#18	CIN#8	1.37722e-17
C791	net6#5	VDD	1.36015e-17
C792	net6	VDD	1.94679e-17
C793	net7#9	PHI#1	1.00222e-18
C794	net8#3	VDD	1.12868e-17
C795	net18#2	VDD#23	1.22651e-18
C796	net1	VDD	2.43487e-17
C797	net3#6	VDD	8.10974e-18
C798	GND#37	COUT	1.81371e-17
C799	net2#20	SOUT#8	4.85966e-17
C800	GND#34	RST#1	4.78312e-19
C801	CIN#4	VDD	1.90404e-17
C802	SOUT#15	VDD#54	1.00955e-16
C803	COUT#12	GND#31	9.33149e-18
C804	COUT#9	net3#4	7.42723e-18
C805	net7	VDD	2.5565e-17
C806	net4#13	VDD#43	1.37551e-17
C807	GND#8	net7#9	1.69099e-18
C808	net10#6	GND#35	7.62312e-17
C809	net13#8	net13#6	1.14012e-18
C810	CIN#10	net3#14	1.36342e-17
C811	net14#12	net3#5	6.93363e-18
C812	net3#7	GND#42	8.05725e-18
C813	net14#11	VDD#37	8.28564e-18
C814	net1#13	net1#3	1.98787e-18
C815	VDD#44	net4#7	2.65072e-18
C816	net1#5	net1	1.68117e-18
C817	VDD#11	net13#8	3.82828e-18
C818	net2#9	net2#10	1.55687e-17
C819	net2#20	net37#6	2.28415e-18
C820	VDD#22	net6	1.63378e-18
C821	net2#8	net2#10	4.86829e-18
C822	RST	VDD	1.14301e-18
C823	net5	net5#3	4.89701e-18
C824	net4#13	VDD#17	2.36805e-17
C825	net2#22	CIN#6	6.53224e-18
C826	VDD#51	net6	3.76291e-18
C827	net6#10	CIN#10	5.61765e-18
C828	VDD#16	net27#8	6.86059e-18
C829	SOUT#15	VDD#3	3.71003e-18
C830	VDD#40	net14#12	2.17431e-17
C831	COUT#9	COUT#8	2.72909e-18
C832	SOUT#15	CIN#3	4.07308e-18
C833	GND#22	GND	1.3387e-17
C834	GND#35	GND	9.10424e-17
C835	net8#9	net8#10	1.28474e-17
C836	GND#16	GND	1.60547e-17
C837	GND#31	GND	2.7127e-17
C838	GND#34	GND	5.88524e-17
C839	net8#9	net8#13	6.02825e-18
C840	net27#5	net4	4.00127e-18
C841	net5#6	net1#11	1.13125e-17
C842	net27#2	VDD	1.73855e-17
C843	GND#9	GND	1.4077e-17
C844	net1#15	net7#3	6.59356e-18
C845	net13#5	SOUT#1	8.35757e-19
C846	net1#13	net1#15	1.51047e-17
C847	net13#6	net13#2	3.35293e-18
C848	VDD#13	net27#5	2.51834e-17
C849	net27#5	PHI#5	7.36087e-19
C850	net27#5	net4#9	4.67955e-17
C851	net1#15	net7#2	1.11997e-17
C852	net13#2	VDD#52	1.34866e-17
C853	net27#5	VDD#43	6.06296e-18
C854	net1#2	net5#6	1.29196e-17
C855	GND#36	GND	8.90971e-17
C856	net27#2	net4	7.78123e-19
C857	GND#42	GND	2.12995e-16
C858	net1#15	net5#8	8.7953e-19
C859	net13#5	VDD#11	5.34371e-19
C860	net13#5	VDD	1.30491e-18
C861	GND#4	GND	2.90693e-17
C862	net5#6	net1	4.3205e-18
C863	net1#15	net5#2	1.47503e-18
C864	VDD#39	net5#2	3.65782e-19
C865	GND#39	GND	5.64861e-17
C866	net5#6	net5#5	1.0726e-17
C867	net7#9	net27#2	1.16334e-17
C868	net1#15	net12#3	5.17242e-17
C869	net8#9	VDD	3.2968e-17
C870	GND#19	GND	1.83306e-17
C871	net13#2	VDD	1.52325e-17
C872	net13#5	net2#20	3.87072e-18
C873	GND#24	GND	1.25687e-16
C874	net13#2	net13#3	1.21238e-17
C875	net5#2	net7	5.65623e-18
C876	net5#6	VDD	1.75573e-17
C877	GND#38	GND	8.88097e-17
C878	net1#10	net27#2	1.02568e-18
C879	VDD#8	net13#5	4.02796e-17
C880	GND#17	GND	2.3656e-17
C881	net27#5	VDD#14	3.29631e-17
C882	net13#5	net13#6	1.32592e-17
C883	net13#5	net13	6.45813e-19
C884	net27#5	VDD#44	5.08885e-18
C885	net27#5	net4#2	1.17455e-18
C886	GND#27	GND	1.12043e-16
C887	net12#5	net1#15	1.38691e-17
C888	net13#5	SOUT#2	9.32097e-19
C889	GND#8	GND	2.4528e-17
C890	net5#2	VDD	2.57085e-17
C891	GND#25	GND	8.74567e-17
C892	net27#2	net27#3	1.55763e-17
C893	net13#5	net13#2	4.48287e-18
C894	VDD#39	net5#6	8.3063e-19
C895	net5#6	net7#2	1.15715e-18
C896	net5#6	VDD#40	1.24682e-18
C897	net4#9	net27#2	6.94565e-18
C898	net27#2	PHI#5	7.33541e-19
C899	GND#37	GND	1.5535e-16
C900	net27#5	PHI#4	4.47776e-19
C901	net27#2	net1#4	8.48232e-18
C902	net5#2	net5#3	1.09952e-17
C903	GND#29	GND	1.80317e-16
C904	net27#2	PHI#4	5.98926e-18
C905	net13#2	net2#19	1.87116e-17
C906	net27#2	VDD#43	2.30456e-17
C907	net5#6	VDD#30	3.1012e-17
C908	GND#1	GND	3.70158e-17
C909	net5#6	net5#9	6.00515e-19
C910	GND#23	GND	1.36672e-16
C911	net8#9	net7	5.39577e-18
C912	SOUT#8	net13#5	1.99012e-18
C913	net5#6	net7	7.70527e-19
C914	net27#5	VDD	1.64755e-17
C915	GND#28	GND	1.45681e-16
C916	net1#11	net5#2	2.86017e-17
C917	net13#5	VDD#53	3.74239e-18
C918	GND#41	GND	9.08373e-17
C919	net5#2	net8#9	5.03196e-17
C920	VDD#29	net5#6	2.47923e-17
C921	net12#3	net8#9	1.53652e-18
C922	net7#9	net27#5	6.45096e-18
C923	GND#11	GND	2.69555e-17
C924	net27#2	net1#5	5.40337e-17
C925	net13#5	net13#9	5.55936e-19
C926	net5#6	net1#9	2.26965e-17
C927	net7#2	net5#2	5.64952e-18
C928	net13#2	SOUT#1	5.78977e-19
C929	net27#5	net27#6	8.38652e-18
C930	net5#2	net1	5.18377e-19
C931	GND#14	GND	7.06671e-18
C932	GND#30	GND	2.96947e-17
C933	net1#9	net5#2	2.5292e-17
C934	GND#5	GND	9.02453e-18
C935	net13#2	net2#9	6.23621e-17
C936	net1#15	net1#14	5.51468e-18
C937	GND#33	GND	2.38504e-17
C938	COUT#13	CIN#4	6.41169e-19
C939	GND#17	CIN#10	1.2376e-18
C940	GND#11	CIN#2	1.48281e-18
C941	VDD#26	CIN#10	1.25566e-18
C942	CIN#8	net2#13	1.0502e-18
C943	net2#18	CIN#5	1.05702e-18
C944	net2#13	CIN#4	1.48154e-18
C945	COUT#4	VDD#33	7.09852e-19
C946	COUT#3	VDD#33	7.2578e-19
C947	COUT#7	VDD#34	7.63515e-19
C948	COUT#7	VDD#37	8.0203e-19
C949	VDD#34	COUT#11	1.09511e-18
C950	VDD#38	COUT#10	1.11577e-18
C951	COUT#4	VDD#40	1.21121e-18
C952	GND#17	SOUT#17	1.0527e-18
C953	GND#35	SOUT#3	1.2522e-18
C954	GND#14	VDD#25	1.07325e-18
C955	GND#5	VDD#11	1.0798e-18
C956	GND#19	VDD#30	1.08184e-18
C957	GND#8	VDD#14	1.11398e-18
C958	GND#8	VDD#16	1.30319e-18
C959	GND#19	VDD#32	1.39733e-18
C960	VDD#34	GND#22	2.136e-18
C961	VDD#17	GND#9	2.18931e-18
C962	GND#1	VDD#1	2.26001e-18
C963	net2#2	GND#35	1.40231e-18
C964	net18#11	CIN#5	1.69058e-19
C965	net18#2	CIN#4	1.89292e-19
C966	net18	CIN#4	3.12001e-19
C967	CIN#8	net18#6	3.23488e-19
C968	VDD#28	PHI#4	4.47088e-19
C969	VDD#13	PHI#2	5.82722e-19
C970	VDD#14	PHI#1	6.24749e-19
C971	VDD#32	PHI#4	7.02357e-19
C972	VDD#13	PHI#1	7.24981e-19
C973	VDD#29	PHI#4	7.80422e-19
C974	COUT#12	net6#5	8.49968e-19
C975	net5#8	net1	3.00311e-19
C976	COUT#10	net3#5	5.05243e-19
C977	COUT#1	net3#4	8.67149e-19
C978	net3#12	COUT#1	9.033e-19
C979	COUT#12	net3#4	1.07146e-18
C980	COUT#4	net3#6	1.28577e-18
C981	VDD#52	SOUT#6	8.44997e-19
C982	VDD#8	SOUT#2	1.18857e-18
C983	VDD#7	SOUT#1	1.36878e-18
C984	VDD#11	SOUT#1	1.54565e-18
C985	SOUT#8	VDD#11	1.7286e-18
C986	net4	PHI#4	4.67721e-19
C987	net4#2	PHI#4	4.73002e-19
C988	GND#22	net6#4	1.25005e-18
C989	net2#19	SOUT#1	6.39923e-19
C990	net2#20	SOUT#3	1.5295e-18
C991	GND#30	net3#4	1.49234e-18
C992	GND#22	net3#5	1.50649e-18
C993	GND#34	net3#3	1.6421e-18
C994	net3#16	GND#14	1.7846e-18
C995	net4#4	RST#2	2.52157e-19
C996	VDD#6	net2#2	7.83973e-19
C997	VDD#8	net2#20	9.14113e-19
C998	VDD#17	net2#3	9.65676e-19
C999	net2#2	VDD	1.3771e-18
C1000	GND#38	net8	2.22149e-18
C1001	net4#9	VDD#16	7.47006e-19
C1002	net6#10	SOUT#6	1.3567e-18
C1003	net27#8	PHI#4	3.12142e-19
C1004	net6#10	VDD#23	8.14423e-19
C1005	net6#10	VDD#21	8.48489e-19
C1006	VDD#40	net6#5	1.16019e-18
C1007	net6#9	VDD#52	1.38283e-18
C1008	SOUT#3	net3#3	5.76547e-19
C1009	VDD#22	net3#16	9.09654e-19
C1010	VDD#20	net3#14	9.78488e-19
C1011	VDD#26	net3#13	9.87129e-19
C1012	VDD#33	net3#6	1.38172e-18
C1013	VDD#37	net3#6	1.49028e-18
C1014	VDD#39	net3#6	1.68758e-18
C1015	VDD#52	net3	1.91607e-18
C1016	net2#22	net6#2	4.48328e-19
C1017	net6#13	net2#7	5.09814e-19
C1018	net6#13	net2#12	8.90317e-19
C1019	net2#7	net6#2	1.02342e-18
C1020	net2#9	net6	1.03882e-18
C1021	net6#10	net2#8	1.2991e-18
C1022	net1#5	net7#2	8.19104e-19
C1023	SOUT#17	net8	9.54038e-19
C1024	SOUT#9	net8#2	1.0179e-18
C1025	net2#14	net18#10	3.37566e-19
C1026	net5#10	net7	3.00311e-19
C1027	net6#13	net3#2	6.42151e-19
C1028	net6#5	net3#5	6.85888e-19
C1029	net6#10	net3	6.96404e-19
C1030	net6#4	net3#4	8.10669e-19
C1031	net6#5	net3#6	8.2065e-19
C1032	net6#13	net3	9.20573e-19
C1033	net3#12	net6#3	1.15477e-18
C1034	net18#7	net6	1.9849e-19
C1035	net6#13	net18#3	2.55286e-19
C1036	net18#2	net6	2.77523e-19
C1037	net18#6	net6	3.22577e-19
C1038	net14#2	net3#12	3.94481e-19
C1039	CIN	GND	4.04619e-17
C1040	COUT	GND	5.04212e-17
C1041	PHI	GND	2.67871e-17
C1042	RST	GND	6.65071e-17
C1043	SOUT	GND	4.66214e-17
C1044	VDD	GND	3.3079e-18
C1045	net7	GND	1.0175e-18
C1046	CIN#4	GND	2.62216e-18
C1047	net3#6	GND	1.6289e-18
C1048	net1	GND	1.34619e-18
C1049	net8#3	GND	2.80962e-18
C1050	net6	GND	5.80245e-18
C1051	net6#5	GND	8.17129e-18
C1052	PHI#4	GND	1.15824e-18
C1053	RST#3	GND	3.14168e-18
C1054	net3	GND	1.13992e-17
C1055	net4	GND	3.12142e-19
C1056	SOUT#1	GND	4.90303e-19
C1057	net2#3	GND	6.98949e-19
C1058	CIN#3	GND	4.78921e-18
C1059	net7#3	GND	1.94396e-17
C1060	CIN#6	GND	1.61542e-17
C1061	net3#4	GND	1.32676e-17
C1062	net1#3	GND	3.51203e-17
C1063	net8	GND	2.0439e-17
C1064	net6#2	GND	4.4656e-17
C1065	net6#4	GND	2.22843e-17
C1066	PHI#6	GND	1.56234e-17
C1067	SOUT#4	GND	2.78191e-17
C1068	RST#1	GND	1.36737e-17
C1069	net3#3	GND	1.56154e-17
C1070	net4#3	GND	2.78771e-17
C1071	SOUT#3	GND	1.33513e-17
C1072	net2	GND	5.04393e-18
C1073	CIN#1	GND	1.76453e-17
C1074	PHI#3	GND	9.84236e-18
C1075	net7#2	GND	1.25313e-16
C1076	CIN#5	GND	3.45253e-17
C1077	net3#5	GND	1.13859e-17
C1078	net1#2	GND	1.2026e-17
C1079	net8#2	GND	7.40327e-17
C1080	net6#3	GND	5.75678e-17
C1081	PHI#5	GND	6.99282e-17
C1082	SOUT#5	GND	2.63043e-17
C1083	RST#2	GND	4.85676e-17
C1084	net3#2	GND	1.89119e-17
C1085	net4#2	GND	1.04124e-17
C1086	SOUT#2	GND	4.32458e-17
C1087	net2#2	GND	2.39851e-17
C1088	CIN#2	GND	1.40695e-16
C1089	PHI#2	GND	8.6089e-17
C1090	VDD#47	GND	1.80586e-17
C1091	VDD#38	GND	1.46911e-17
C1092	net8#6	GND	8.65059e-17
C1093	net8#13	GND	3.90235e-17
C1094	net8#14	GND	1.73409e-16
C1095	COUT#10	GND	1.57504e-16
C1096	COUT#13	GND	4.7741e-17
C1097	net3#13	GND	1.15356e-16
C1098	net3#15	GND	3.2808e-17
C1099	net12#3	GND	5.90619e-18
C1100	net12#5	GND	7.47594e-17
C1101	net8#9	GND	6.04217e-19
C1102	CIN#10	GND	5.45319e-17
C1103	CIN#8	GND	2.94989e-17
C1104	net1#9	GND	3.08046e-18
C1105	net1#11	GND	4.4866e-18
C1106	net1#13	GND	1.45404e-17
C1107	net2#18	GND	1.81906e-18
C1108	net2#22	GND	2.03996e-17
C1109	net2#14	GND	1.558e-18
C1110	COUT#9	GND	1.66341e-17
C1111	COUT#11	GND	5.33636e-17
C1112	net14#9	GND	5.18511e-20
C1113	net14#11	GND	5.01504e-19
C1114	net18#11	GND	1.77714e-18
C1115	net18#7	GND	9.71176e-19
C1116	net37#4	GND	1.26365e-17
C1117	net37#5	GND	6.43795e-17
C1118	VDD#34	GND	9.1376e-19
C1119	VDD#39	GND	6.41572e-20
C1120	SOUT#17	GND	1.83378e-17
C1121	SOUT#13	GND	1.92132e-18
C1122	net21#3	GND	1.41957e-17
C1123	net21#5	GND	2.3838e-17
C1124	SOUT#9	GND	1.28794e-17
C1125	SOUT#11	GND	4.01254e-18
C1126	SOUT#14	GND	3.79279e-18
C1127	VDD#40	GND	1.87382e-19
C1128	VDD#29	GND	8.06149e-19
C1129	VDD#50	GND	8.39147e-19
C1130	COUT#4	GND	9.14475e-19
C1131	net18#12	GND	2.91229e-18
C1132	net18#2	GND	3.0103e-18
C1133	net33#5	GND	3.03995e-17
C1134	net33#3	GND	5.05107e-18
C1135	COUT#1	GND	7.49483e-18
C1136	COUT#12	GND	2.46811e-17
C1137	VDD#22	GND	1.65055e-18
C1138	net14#2	GND	3.18649e-18
C1139	net14#12	GND	1.7817e-18
C1140	net6#10	GND	2.44372e-17
C1141	net6#13	GND	4.15562e-17
C1142	net3#16	GND	4.87025e-17
C1143	net3#12	GND	2.32379e-17
C1144	net1#10	GND	2.16671e-18
C1145	net1#5	GND	1.49748e-19
C1146	net21	GND	1.99362e-17
C1147	net21#6	GND	2.54695e-17
C1148	net6#7	GND	2.06191e-17
C1149	net6#11	GND	1.51734e-17
C1150	net27#2	GND	1.81345e-18
C1151	net8#4	GND	2.01708e-17
C1152	net8#15	GND	5.65615e-17
C1153	net10#5	GND	2.92884e-17
C1154	net10#3	GND	6.14473e-18
C1155	net4#12	GND	5.39045e-18
C1156	net4#11	GND	1.54664e-18
C1157	net2#9	GND	3.14112e-19
C1158	VDD#52	GND	5.40178e-19
C1159	net2#19	GND	5.401e-18
C1160	net2#7	GND	6.62161e-18
C1161	net13#2	GND	7.57215e-18
C1162	net33#6	GND	2.99855e-17
C1163	net33	GND	1.15404e-17
C1164	net4#13	GND	6.98949e-19
C1165	net4#9	GND	2.92698e-18
C1166	net27#5	GND	2.07877e-18
C1167	net12#2	GND	1.87723e-17
C1168	net12#6	GND	7.473e-17
C1169	VDD#13	GND	1.72134e-18
C1170	net13#5	GND	3.86761e-18
C1171	net37#2	GND	1.95679e-17
C1172	net37#6	GND	8.01368e-17
C1173	net4#4	GND	1.47938e-17
C1174	net4#14	GND	3.11895e-18
C1175	net3#7	GND	1.70551e-17
C1176	net3#14	GND	7.74513e-17
C1177	net3#9	GND	7.34082e-18
C1178	VDD#53	GND	5.90251e-19
C1179	VDD#8	GND	6.41686e-19
C1180	net10#6	GND	3.09339e-17
C1181	net10	GND	6.61111e-18
C1182	VDD#6	GND	2.12686e-18
C1183	VDD#54	GND	2.24582e-17
C1184	net2#20	GND	3.035e-17
C1185	net2#5	GND	5.05974e-17
C1186	SOUT#8	GND	4.52341e-17
C1187	SOUT#15	GND	3.84121e-19
C1188	net7#9	GND	8.00536e-17
C1189	net7#5	GND	5.95288e-19
C1190	net7#6	GND	1.72011e-17
C1191	VDD#46	GND	2.12717e-17
C1192	net8#10	GND	5.90088e-19
C1193	net2#15	GND	6.11864e-19
C1194	net14#7	GND	1.01697e-19
C1195	net18#8	GND	3.47442e-19
C1196	VDD#35	GND	2.13299e-19
C1197	net5#5	GND	1.43426e-19
C1198	COUT#5	GND	2.95659e-22
C1199	VDD#23	GND	8.26354e-19
C1200	net14#3	GND	1.33231e-18
C1201	net27#3	GND	4.77501e-19
C1202	net13#3	GND	2.14104e-20
C1203	net27#6	GND	1.32517e-19
C1204	VDD#14	GND	1.15206e-19
C1205	net13#6	GND	1.56041e-18
C1206	VDD#9	GND	2.75182e-19
C1207	net21#4	GND	1.7731e-19
C1208	net33#2	GND	4.75427e-20
C1209	net12	GND	3.66612e-20
C1210	net37	GND	2.39008e-19
C1211	VDD#11	GND	6.49289e-20
C1212	VDD#7	GND	1.26994e-18
C1213	VDD#12	GND	4.62384e-19
C1214	net13#8	GND	1.43177e-18
C1215	net13#9	GND	2.6831e-18
C1216	net13	GND	1.91584e-18
C1217	net2#12	GND	3.12901e-19
C1218	net2#8	GND	2.95349e-19
C1219	net27#8	GND	7.80348e-19
C1220	net27#9	GND	2.51134e-19
C1221	net27	GND	1.39967e-18
C1222	net1#8	GND	2.27423e-19
C1223	net1#4	GND	2.6882e-20
C1224	VDD#25	GND	3.39718e-19
C1225	VDD#21	GND	2.48665e-19
C1226	net14#5	GND	4.31334e-19
C1227	net14	GND	1.50953e-18
C1228	net18#5	GND	1.07806e-18
C1229	COUT#7	GND	3.48418e-19
C1230	COUT#3	GND	4.22926e-19
C1231	VDD#37	GND	4.54904e-19
C1232	VDD#33	GND	9.24701e-19
C1233	SOUT#16	GND	1.75015e-18
C1234	net18#10	GND	8.84065e-19
C1235	net14#10	GND	6.75463e-20
C1236	net14#6	GND	8.64449e-20
C1237	net2#17	GND	1.12478e-18
C1238	net2#13	GND	1.99284e-19
C1239	net5#9	GND	7.40201e-19
C1240	net5	GND	2.54561e-19
C1241	net5#6	GND	2.60389e-18
C1242	net1#15	GND	1.34079e-17
C1243	net8#12	GND	6.47031e-19
C1244	net8#8	GND	5.95537e-19
*
*
.ENDS XOR_X1
*
